// unnamed.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module unnamed (
		output wire [13:0]  araddr,   // altera_axi4_master.araddr
		output wire [1:0]   arburst,  //                   .arburst
		output wire [3:0]   arcache,  //                   .arcache
		output wire         arid,     //                   .arid
		output wire [7:0]   arlen,    //                   .arlen
		output wire         arlock,   //                   .arlock
		output wire [2:0]   arprot,   //                   .arprot
		output wire [3:0]   arqos,    //                   .arqos
		input  wire         arready,  //                   .arready
		output wire [3:0]   arregion, //                   .arregion
		output wire [2:0]   arsize,   //                   .arsize
		output wire         arvalid,  //                   .arvalid
		output wire [13:0]  awaddr,   //                   .awaddr
		output wire [1:0]   awburst,  //                   .awburst
		output wire [3:0]   awcache,  //                   .awcache
		output wire         awid,     //                   .awid
		output wire [7:0]   awlen,    //                   .awlen
		output wire         awlock,   //                   .awlock
		output wire [2:0]   awprot,   //                   .awprot
		output wire [3:0]   awqos,    //                   .awqos
		input  wire         awready,  //                   .awready
		output wire [3:0]   awregion, //                   .awregion
		output wire [2:0]   awsize,   //                   .awsize
		output wire         awvalid,  //                   .awvalid
		input  wire         bid,      //                   .bid
		output wire         bready,   //                   .bready
		input  wire [1:0]   bresp,    //                   .bresp
		input  wire         bvalid,   //                   .bvalid
		input  wire [127:0] rdata,    //                   .rdata
		input  wire         rid,      //                   .rid
		input  wire         rlast,    //                   .rlast
		output wire         rready,   //                   .rready
		input  wire [1:0]   rresp,    //                   .rresp
		input  wire         rvalid,   //                   .rvalid
		output wire [127:0] wdata,    //                   .wdata
		output wire         wlast,    //                   .wlast
		input  wire         wready,   //                   .wready
		output wire [15:0]  wstrb,    //                   .wstrb
		output wire         wvalid,   //                   .wvalid
		input  wire         CLK,      //              clock.clk
		input  wire         RST_N     //         reset_sink.reset_n
	);

	unnamed_axiMaster_0 aximaster_0 (
		.CLK      (CLK),      //              clock.clk
		.araddr   (araddr),   // altera_axi4_master.araddr
		.arburst  (arburst),  //                   .arburst
		.arcache  (arcache),  //                   .arcache
		.arid     (arid),     //                   .arid
		.arlen    (arlen),    //                   .arlen
		.arlock   (arlock),   //                   .arlock
		.arprot   (arprot),   //                   .arprot
		.arqos    (arqos),    //                   .arqos
		.arready  (arready),  //                   .arready
		.arregion (arregion), //                   .arregion
		.arsize   (arsize),   //                   .arsize
		.arvalid  (arvalid),  //                   .arvalid
		.awaddr   (awaddr),   //                   .awaddr
		.awburst  (awburst),  //                   .awburst
		.awcache  (awcache),  //                   .awcache
		.awid     (awid),     //                   .awid
		.awlen    (awlen),    //                   .awlen
		.awlock   (awlock),   //                   .awlock
		.awprot   (awprot),   //                   .awprot
		.awqos    (awqos),    //                   .awqos
		.awready  (awready),  //                   .awready
		.awregion (awregion), //                   .awregion
		.awsize   (awsize),   //                   .awsize
		.awvalid  (awvalid),  //                   .awvalid
		.bid      (bid),      //                   .bid
		.bready   (bready),   //                   .bready
		.bresp    (bresp),    //                   .bresp
		.bvalid   (bvalid),   //                   .bvalid
		.rdata    (rdata),    //                   .rdata
		.rid      (rid),      //                   .rid
		.rlast    (rlast),    //                   .rlast
		.rready   (rready),   //                   .rready
		.rresp    (rresp),    //                   .rresp
		.rvalid   (rvalid),   //                   .rvalid
		.wdata    (wdata),    //                   .wdata
		.wlast    (wlast),    //                   .wlast
		.wready   (wready),   //                   .wready
		.wstrb    (wstrb),    //                   .wstrb
		.wvalid   (wvalid),   //                   .wvalid
		.RST_N    (RST_N)     //         reset_sink.reset_n
	);

endmodule
