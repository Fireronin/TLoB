
module Example1B (
	clk_clk,
	reset_reset_n,
	simplefifo_2_enq_en_wire);	

	input		clk_clk;
	input		reset_reset_n;
	input		simplefifo_2_enq_en_wire;
endmodule
