-- Example3.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Example3 is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity Example3;

architecture rtl of Example3 is
	component Example3_axi4Slave_0 is
		port (
			CLK      : in  std_logic                      := 'X';             -- clk
			araddr   : in  std_logic_vector(13 downto 0)  := (others => 'X'); -- araddr
			arburst  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			arcache  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			arid     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arid
			arlen    : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- arlen
			arlock   : in  std_logic                      := 'X';             -- arlock
			arprot   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			arqos    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arqos
			arready  : out std_logic;                                         -- arready
			arregion : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arregion
			arsize   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			arvalid  : in  std_logic                      := 'X';             -- arvalid
			awaddr   : in  std_logic_vector(13 downto 0)  := (others => 'X'); -- awaddr
			awburst  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			awcache  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			awid     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awid
			awlen    : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- awlen
			awlock   : in  std_logic                      := 'X';             -- awlock
			awprot   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			awqos    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awqos
			awready  : out std_logic;                                         -- awready
			awregion : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awregion
			awsize   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			awvalid  : in  std_logic                      := 'X';             -- awvalid
			bid      : out std_logic_vector(1 downto 0);                      -- bid
			bready   : in  std_logic                      := 'X';             -- bready
			bresp    : out std_logic_vector(1 downto 0);                      -- bresp
			bvalid   : out std_logic;                                         -- bvalid
			rdata    : out std_logic_vector(127 downto 0);                    -- rdata
			rid      : out std_logic_vector(1 downto 0);                      -- rid
			rlast    : out std_logic;                                         -- rlast
			rready   : in  std_logic                      := 'X';             -- rready
			rresp    : out std_logic_vector(1 downto 0);                      -- rresp
			rvalid   : out std_logic;                                         -- rvalid
			wdata    : in  std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			wlast    : in  std_logic                      := 'X';             -- wlast
			wready   : out std_logic;                                         -- wready
			wstrb    : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			wvalid   : in  std_logic                      := 'X';             -- wvalid
			RST_N    : in  std_logic                      := 'X'              -- reset_n
		);
	end component Example3_axi4Slave_0;

	component Example3_axiMaster_0 is
		port (
			CLK      : in  std_logic                      := 'X';             -- clk
			araddr   : out std_logic_vector(13 downto 0);                     -- araddr
			arburst  : out std_logic_vector(1 downto 0);                      -- arburst
			arcache  : out std_logic_vector(3 downto 0);                      -- arcache
			arid     : out std_logic;                                         -- arid
			arlen    : out std_logic_vector(7 downto 0);                      -- arlen
			arlock   : out std_logic;                                         -- arlock
			arprot   : out std_logic_vector(2 downto 0);                      -- arprot
			arqos    : out std_logic_vector(3 downto 0);                      -- arqos
			arready  : in  std_logic                      := 'X';             -- arready
			arregion : out std_logic_vector(3 downto 0);                      -- arregion
			arsize   : out std_logic_vector(2 downto 0);                      -- arsize
			arvalid  : out std_logic;                                         -- arvalid
			awaddr   : out std_logic_vector(13 downto 0);                     -- awaddr
			awburst  : out std_logic_vector(1 downto 0);                      -- awburst
			awcache  : out std_logic_vector(3 downto 0);                      -- awcache
			awid     : out std_logic;                                         -- awid
			awlen    : out std_logic_vector(7 downto 0);                      -- awlen
			awlock   : out std_logic;                                         -- awlock
			awprot   : out std_logic_vector(2 downto 0);                      -- awprot
			awqos    : out std_logic_vector(3 downto 0);                      -- awqos
			awready  : in  std_logic                      := 'X';             -- awready
			awregion : out std_logic_vector(3 downto 0);                      -- awregion
			awsize   : out std_logic_vector(2 downto 0);                      -- awsize
			awvalid  : out std_logic;                                         -- awvalid
			bid      : in  std_logic                      := 'X';             -- bid
			bready   : out std_logic;                                         -- bready
			bresp    : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			bvalid   : in  std_logic                      := 'X';             -- bvalid
			rdata    : in  std_logic_vector(127 downto 0) := (others => 'X'); -- rdata
			rid      : in  std_logic                      := 'X';             -- rid
			rlast    : in  std_logic                      := 'X';             -- rlast
			rready   : out std_logic;                                         -- rready
			rresp    : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			rvalid   : in  std_logic                      := 'X';             -- rvalid
			wdata    : out std_logic_vector(127 downto 0);                    -- wdata
			wlast    : out std_logic;                                         -- wlast
			wready   : in  std_logic                      := 'X';             -- wready
			wstrb    : out std_logic_vector(15 downto 0);                     -- wstrb
			wvalid   : out std_logic;                                         -- wvalid
			RST_N    : in  std_logic                      := 'X'              -- reset_n
		);
	end component Example3_axiMaster_0;

	component Example3_mm_interconnect_0 is
		port (
			axi4Slave_0_altera_axi4_slave_awid                 : out std_logic_vector(1 downto 0);                      -- awid
			axi4Slave_0_altera_axi4_slave_awaddr               : out std_logic_vector(13 downto 0);                     -- awaddr
			axi4Slave_0_altera_axi4_slave_awlen                : out std_logic_vector(7 downto 0);                      -- awlen
			axi4Slave_0_altera_axi4_slave_awsize               : out std_logic_vector(2 downto 0);                      -- awsize
			axi4Slave_0_altera_axi4_slave_awburst              : out std_logic_vector(1 downto 0);                      -- awburst
			axi4Slave_0_altera_axi4_slave_awlock               : out std_logic_vector(0 downto 0);                      -- awlock
			axi4Slave_0_altera_axi4_slave_awcache              : out std_logic_vector(3 downto 0);                      -- awcache
			axi4Slave_0_altera_axi4_slave_awprot               : out std_logic_vector(2 downto 0);                      -- awprot
			axi4Slave_0_altera_axi4_slave_awqos                : out std_logic_vector(3 downto 0);                      -- awqos
			axi4Slave_0_altera_axi4_slave_awregion             : out std_logic_vector(3 downto 0);                      -- awregion
			axi4Slave_0_altera_axi4_slave_awvalid              : out std_logic;                                         -- awvalid
			axi4Slave_0_altera_axi4_slave_awready              : in  std_logic                      := 'X';             -- awready
			axi4Slave_0_altera_axi4_slave_wdata                : out std_logic_vector(127 downto 0);                    -- wdata
			axi4Slave_0_altera_axi4_slave_wstrb                : out std_logic_vector(15 downto 0);                     -- wstrb
			axi4Slave_0_altera_axi4_slave_wlast                : out std_logic;                                         -- wlast
			axi4Slave_0_altera_axi4_slave_wvalid               : out std_logic;                                         -- wvalid
			axi4Slave_0_altera_axi4_slave_wready               : in  std_logic                      := 'X';             -- wready
			axi4Slave_0_altera_axi4_slave_bid                  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- bid
			axi4Slave_0_altera_axi4_slave_bresp                : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			axi4Slave_0_altera_axi4_slave_bvalid               : in  std_logic                      := 'X';             -- bvalid
			axi4Slave_0_altera_axi4_slave_bready               : out std_logic;                                         -- bready
			axi4Slave_0_altera_axi4_slave_arid                 : out std_logic_vector(1 downto 0);                      -- arid
			axi4Slave_0_altera_axi4_slave_araddr               : out std_logic_vector(13 downto 0);                     -- araddr
			axi4Slave_0_altera_axi4_slave_arlen                : out std_logic_vector(7 downto 0);                      -- arlen
			axi4Slave_0_altera_axi4_slave_arsize               : out std_logic_vector(2 downto 0);                      -- arsize
			axi4Slave_0_altera_axi4_slave_arburst              : out std_logic_vector(1 downto 0);                      -- arburst
			axi4Slave_0_altera_axi4_slave_arlock               : out std_logic_vector(0 downto 0);                      -- arlock
			axi4Slave_0_altera_axi4_slave_arcache              : out std_logic_vector(3 downto 0);                      -- arcache
			axi4Slave_0_altera_axi4_slave_arprot               : out std_logic_vector(2 downto 0);                      -- arprot
			axi4Slave_0_altera_axi4_slave_arqos                : out std_logic_vector(3 downto 0);                      -- arqos
			axi4Slave_0_altera_axi4_slave_arregion             : out std_logic_vector(3 downto 0);                      -- arregion
			axi4Slave_0_altera_axi4_slave_arvalid              : out std_logic;                                         -- arvalid
			axi4Slave_0_altera_axi4_slave_arready              : in  std_logic                      := 'X';             -- arready
			axi4Slave_0_altera_axi4_slave_rid                  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rid
			axi4Slave_0_altera_axi4_slave_rdata                : in  std_logic_vector(127 downto 0) := (others => 'X'); -- rdata
			axi4Slave_0_altera_axi4_slave_rresp                : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			axi4Slave_0_altera_axi4_slave_rlast                : in  std_logic                      := 'X';             -- rlast
			axi4Slave_0_altera_axi4_slave_rvalid               : in  std_logic                      := 'X';             -- rvalid
			axi4Slave_0_altera_axi4_slave_rready               : out std_logic;                                         -- rready
			axiMaster_0_altera_axi4_master_awid                : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- awid
			axiMaster_0_altera_axi4_master_awaddr              : in  std_logic_vector(13 downto 0)  := (others => 'X'); -- awaddr
			axiMaster_0_altera_axi4_master_awlen               : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- awlen
			axiMaster_0_altera_axi4_master_awsize              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			axiMaster_0_altera_axi4_master_awburst             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			axiMaster_0_altera_axi4_master_awlock              : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- awlock
			axiMaster_0_altera_axi4_master_awcache             : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			axiMaster_0_altera_axi4_master_awprot              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			axiMaster_0_altera_axi4_master_awqos               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awqos
			axiMaster_0_altera_axi4_master_awregion            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awregion
			axiMaster_0_altera_axi4_master_awvalid             : in  std_logic                      := 'X';             -- awvalid
			axiMaster_0_altera_axi4_master_awready             : out std_logic;                                         -- awready
			axiMaster_0_altera_axi4_master_wdata               : in  std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			axiMaster_0_altera_axi4_master_wstrb               : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			axiMaster_0_altera_axi4_master_wlast               : in  std_logic                      := 'X';             -- wlast
			axiMaster_0_altera_axi4_master_wvalid              : in  std_logic                      := 'X';             -- wvalid
			axiMaster_0_altera_axi4_master_wready              : out std_logic;                                         -- wready
			axiMaster_0_altera_axi4_master_bid                 : out std_logic_vector(0 downto 0);                      -- bid
			axiMaster_0_altera_axi4_master_bresp               : out std_logic_vector(1 downto 0);                      -- bresp
			axiMaster_0_altera_axi4_master_bvalid              : out std_logic;                                         -- bvalid
			axiMaster_0_altera_axi4_master_bready              : in  std_logic                      := 'X';             -- bready
			axiMaster_0_altera_axi4_master_arid                : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- arid
			axiMaster_0_altera_axi4_master_araddr              : in  std_logic_vector(13 downto 0)  := (others => 'X'); -- araddr
			axiMaster_0_altera_axi4_master_arlen               : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- arlen
			axiMaster_0_altera_axi4_master_arsize              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			axiMaster_0_altera_axi4_master_arburst             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			axiMaster_0_altera_axi4_master_arlock              : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- arlock
			axiMaster_0_altera_axi4_master_arcache             : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			axiMaster_0_altera_axi4_master_arprot              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			axiMaster_0_altera_axi4_master_arqos               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arqos
			axiMaster_0_altera_axi4_master_arregion            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arregion
			axiMaster_0_altera_axi4_master_arvalid             : in  std_logic                      := 'X';             -- arvalid
			axiMaster_0_altera_axi4_master_arready             : out std_logic;                                         -- arready
			axiMaster_0_altera_axi4_master_rid                 : out std_logic_vector(0 downto 0);                      -- rid
			axiMaster_0_altera_axi4_master_rdata               : out std_logic_vector(127 downto 0);                    -- rdata
			axiMaster_0_altera_axi4_master_rresp               : out std_logic_vector(1 downto 0);                      -- rresp
			axiMaster_0_altera_axi4_master_rlast               : out std_logic;                                         -- rlast
			axiMaster_0_altera_axi4_master_rvalid              : out std_logic;                                         -- rvalid
			axiMaster_0_altera_axi4_master_rready              : in  std_logic                      := 'X';             -- rready
			clk_0_clk_clk                                      : in  std_logic                      := 'X';             -- clk
			axiMaster_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X'              -- reset
		);
	end component Example3_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal aximaster_0_altera_axi4_master_awburst                   : std_logic_vector(1 downto 0);   -- axiMaster_0:awburst -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awburst
	signal aximaster_0_altera_axi4_master_arregion                  : std_logic_vector(3 downto 0);   -- axiMaster_0:arregion -> mm_interconnect_0:axiMaster_0_altera_axi4_master_arregion
	signal aximaster_0_altera_axi4_master_arlen                     : std_logic_vector(7 downto 0);   -- axiMaster_0:arlen -> mm_interconnect_0:axiMaster_0_altera_axi4_master_arlen
	signal aximaster_0_altera_axi4_master_arqos                     : std_logic_vector(3 downto 0);   -- axiMaster_0:arqos -> mm_interconnect_0:axiMaster_0_altera_axi4_master_arqos
	signal aximaster_0_altera_axi4_master_wready                    : std_logic;                      -- mm_interconnect_0:axiMaster_0_altera_axi4_master_wready -> axiMaster_0:wready
	signal aximaster_0_altera_axi4_master_wstrb                     : std_logic_vector(15 downto 0);  -- axiMaster_0:wstrb -> mm_interconnect_0:axiMaster_0_altera_axi4_master_wstrb
	signal aximaster_0_altera_axi4_master_rid                       : std_logic;                      -- mm_interconnect_0:axiMaster_0_altera_axi4_master_rid -> axiMaster_0:rid
	signal aximaster_0_altera_axi4_master_rready                    : std_logic;                      -- axiMaster_0:rready -> mm_interconnect_0:axiMaster_0_altera_axi4_master_rready
	signal aximaster_0_altera_axi4_master_awlen                     : std_logic_vector(7 downto 0);   -- axiMaster_0:awlen -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awlen
	signal aximaster_0_altera_axi4_master_awqos                     : std_logic_vector(3 downto 0);   -- axiMaster_0:awqos -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awqos
	signal aximaster_0_altera_axi4_master_arcache                   : std_logic_vector(3 downto 0);   -- axiMaster_0:arcache -> mm_interconnect_0:axiMaster_0_altera_axi4_master_arcache
	signal aximaster_0_altera_axi4_master_araddr                    : std_logic_vector(13 downto 0);  -- axiMaster_0:araddr -> mm_interconnect_0:axiMaster_0_altera_axi4_master_araddr
	signal aximaster_0_altera_axi4_master_wvalid                    : std_logic;                      -- axiMaster_0:wvalid -> mm_interconnect_0:axiMaster_0_altera_axi4_master_wvalid
	signal aximaster_0_altera_axi4_master_arprot                    : std_logic_vector(2 downto 0);   -- axiMaster_0:arprot -> mm_interconnect_0:axiMaster_0_altera_axi4_master_arprot
	signal aximaster_0_altera_axi4_master_arvalid                   : std_logic;                      -- axiMaster_0:arvalid -> mm_interconnect_0:axiMaster_0_altera_axi4_master_arvalid
	signal aximaster_0_altera_axi4_master_awprot                    : std_logic_vector(2 downto 0);   -- axiMaster_0:awprot -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awprot
	signal aximaster_0_altera_axi4_master_wdata                     : std_logic_vector(127 downto 0); -- axiMaster_0:wdata -> mm_interconnect_0:axiMaster_0_altera_axi4_master_wdata
	signal aximaster_0_altera_axi4_master_arid                      : std_logic;                      -- axiMaster_0:arid -> mm_interconnect_0:axiMaster_0_altera_axi4_master_arid
	signal aximaster_0_altera_axi4_master_awcache                   : std_logic_vector(3 downto 0);   -- axiMaster_0:awcache -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awcache
	signal aximaster_0_altera_axi4_master_arlock                    : std_logic;                      -- axiMaster_0:arlock -> mm_interconnect_0:axiMaster_0_altera_axi4_master_arlock
	signal aximaster_0_altera_axi4_master_awlock                    : std_logic;                      -- axiMaster_0:awlock -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awlock
	signal aximaster_0_altera_axi4_master_awaddr                    : std_logic_vector(13 downto 0);  -- axiMaster_0:awaddr -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awaddr
	signal aximaster_0_altera_axi4_master_arready                   : std_logic;                      -- mm_interconnect_0:axiMaster_0_altera_axi4_master_arready -> axiMaster_0:arready
	signal aximaster_0_altera_axi4_master_bresp                     : std_logic_vector(1 downto 0);   -- mm_interconnect_0:axiMaster_0_altera_axi4_master_bresp -> axiMaster_0:bresp
	signal aximaster_0_altera_axi4_master_rdata                     : std_logic_vector(127 downto 0); -- mm_interconnect_0:axiMaster_0_altera_axi4_master_rdata -> axiMaster_0:rdata
	signal aximaster_0_altera_axi4_master_arburst                   : std_logic_vector(1 downto 0);   -- axiMaster_0:arburst -> mm_interconnect_0:axiMaster_0_altera_axi4_master_arburst
	signal aximaster_0_altera_axi4_master_awready                   : std_logic;                      -- mm_interconnect_0:axiMaster_0_altera_axi4_master_awready -> axiMaster_0:awready
	signal aximaster_0_altera_axi4_master_arsize                    : std_logic_vector(2 downto 0);   -- axiMaster_0:arsize -> mm_interconnect_0:axiMaster_0_altera_axi4_master_arsize
	signal aximaster_0_altera_axi4_master_bready                    : std_logic;                      -- axiMaster_0:bready -> mm_interconnect_0:axiMaster_0_altera_axi4_master_bready
	signal aximaster_0_altera_axi4_master_rlast                     : std_logic;                      -- mm_interconnect_0:axiMaster_0_altera_axi4_master_rlast -> axiMaster_0:rlast
	signal aximaster_0_altera_axi4_master_wlast                     : std_logic;                      -- axiMaster_0:wlast -> mm_interconnect_0:axiMaster_0_altera_axi4_master_wlast
	signal aximaster_0_altera_axi4_master_awregion                  : std_logic_vector(3 downto 0);   -- axiMaster_0:awregion -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awregion
	signal aximaster_0_altera_axi4_master_rresp                     : std_logic_vector(1 downto 0);   -- mm_interconnect_0:axiMaster_0_altera_axi4_master_rresp -> axiMaster_0:rresp
	signal aximaster_0_altera_axi4_master_awid                      : std_logic;                      -- axiMaster_0:awid -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awid
	signal aximaster_0_altera_axi4_master_bid                       : std_logic;                      -- mm_interconnect_0:axiMaster_0_altera_axi4_master_bid -> axiMaster_0:bid
	signal aximaster_0_altera_axi4_master_bvalid                    : std_logic;                      -- mm_interconnect_0:axiMaster_0_altera_axi4_master_bvalid -> axiMaster_0:bvalid
	signal aximaster_0_altera_axi4_master_awsize                    : std_logic_vector(2 downto 0);   -- axiMaster_0:awsize -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awsize
	signal aximaster_0_altera_axi4_master_awvalid                   : std_logic;                      -- axiMaster_0:awvalid -> mm_interconnect_0:axiMaster_0_altera_axi4_master_awvalid
	signal aximaster_0_altera_axi4_master_rvalid                    : std_logic;                      -- mm_interconnect_0:axiMaster_0_altera_axi4_master_rvalid -> axiMaster_0:rvalid
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awburst  : std_logic_vector(1 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awburst -> axi4Slave_0:awburst
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arregion : std_logic_vector(3 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arregion -> axi4Slave_0:arregion
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arlen    : std_logic_vector(7 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arlen -> axi4Slave_0:arlen
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arqos    : std_logic_vector(3 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arqos -> axi4Slave_0:arqos
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_wstrb    : std_logic_vector(15 downto 0);  -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_wstrb -> axi4Slave_0:wstrb
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_wready   : std_logic;                      -- axi4Slave_0:wready -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_wready
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_rid      : std_logic_vector(1 downto 0);   -- axi4Slave_0:rid -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_rid
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_rready   : std_logic;                      -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_rready -> axi4Slave_0:rready
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awlen    : std_logic_vector(7 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awlen -> axi4Slave_0:awlen
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awqos    : std_logic_vector(3 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awqos -> axi4Slave_0:awqos
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arcache  : std_logic_vector(3 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arcache -> axi4Slave_0:arcache
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_wvalid   : std_logic;                      -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_wvalid -> axi4Slave_0:wvalid
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_araddr   : std_logic_vector(13 downto 0);  -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_araddr -> axi4Slave_0:araddr
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arprot   : std_logic_vector(2 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arprot -> axi4Slave_0:arprot
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awprot   : std_logic_vector(2 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awprot -> axi4Slave_0:awprot
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_wdata    : std_logic_vector(127 downto 0); -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_wdata -> axi4Slave_0:wdata
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arvalid  : std_logic;                      -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arvalid -> axi4Slave_0:arvalid
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awcache  : std_logic_vector(3 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awcache -> axi4Slave_0:awcache
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arid     : std_logic_vector(1 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arid -> axi4Slave_0:arid
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arlock   : std_logic_vector(0 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arlock -> axi4Slave_0:arlock
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awlock   : std_logic_vector(0 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awlock -> axi4Slave_0:awlock
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awaddr   : std_logic_vector(13 downto 0);  -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awaddr -> axi4Slave_0:awaddr
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_bresp    : std_logic_vector(1 downto 0);   -- axi4Slave_0:bresp -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_bresp
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arready  : std_logic;                      -- axi4Slave_0:arready -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arready
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_rdata    : std_logic_vector(127 downto 0); -- axi4Slave_0:rdata -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_rdata
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awready  : std_logic;                      -- axi4Slave_0:awready -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awready
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arburst  : std_logic_vector(1 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arburst -> axi4Slave_0:arburst
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_arsize   : std_logic_vector(2 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_arsize -> axi4Slave_0:arsize
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_bready   : std_logic;                      -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_bready -> axi4Slave_0:bready
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_rlast    : std_logic;                      -- axi4Slave_0:rlast -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_rlast
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_wlast    : std_logic;                      -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_wlast -> axi4Slave_0:wlast
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awregion : std_logic_vector(3 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awregion -> axi4Slave_0:awregion
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_rresp    : std_logic_vector(1 downto 0);   -- axi4Slave_0:rresp -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_rresp
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awid     : std_logic_vector(1 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awid -> axi4Slave_0:awid
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_bid      : std_logic_vector(1 downto 0);   -- axi4Slave_0:bid -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_bid
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_bvalid   : std_logic;                      -- axi4Slave_0:bvalid -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_bvalid
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awsize   : std_logic_vector(2 downto 0);   -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awsize -> axi4Slave_0:awsize
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_awvalid  : std_logic;                      -- mm_interconnect_0:axi4Slave_0_altera_axi4_slave_awvalid -> axi4Slave_0:awvalid
	signal mm_interconnect_0_axi4slave_0_altera_axi4_slave_rvalid   : std_logic;                      -- axi4Slave_0:rvalid -> mm_interconnect_0:axi4Slave_0_altera_axi4_slave_rvalid
	signal rst_controller_reset_out_reset                           : std_logic;                      -- rst_controller:reset_out -> [mm_interconnect_0:axiMaster_0_reset_sink_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                  : std_logic;                      -- reset_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv                 : std_logic;                      -- rst_controller_reset_out_reset:inv -> [axi4Slave_0:RST_N, axiMaster_0:RST_N]

begin

	axi4slave_0 : component Example3_axi4Slave_0
		port map (
			CLK      => clk_clk,                                                   --             clock.clk
			araddr   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_araddr,    -- altera_axi4_slave.araddr
			arburst  => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arburst,   --                  .arburst
			arcache  => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arcache,   --                  .arcache
			arid     => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arid,      --                  .arid
			arlen    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arlen,     --                  .arlen
			arlock   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arlock(0), --                  .arlock
			arprot   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arprot,    --                  .arprot
			arqos    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arqos,     --                  .arqos
			arready  => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arready,   --                  .arready
			arregion => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arregion,  --                  .arregion
			arsize   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arsize,    --                  .arsize
			arvalid  => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arvalid,   --                  .arvalid
			awaddr   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awaddr,    --                  .awaddr
			awburst  => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awburst,   --                  .awburst
			awcache  => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awcache,   --                  .awcache
			awid     => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awid,      --                  .awid
			awlen    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awlen,     --                  .awlen
			awlock   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awlock(0), --                  .awlock
			awprot   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awprot,    --                  .awprot
			awqos    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awqos,     --                  .awqos
			awready  => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awready,   --                  .awready
			awregion => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awregion,  --                  .awregion
			awsize   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awsize,    --                  .awsize
			awvalid  => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awvalid,   --                  .awvalid
			bid      => mm_interconnect_0_axi4slave_0_altera_axi4_slave_bid,       --                  .bid
			bready   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_bready,    --                  .bready
			bresp    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_bresp,     --                  .bresp
			bvalid   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_bvalid,    --                  .bvalid
			rdata    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rdata,     --                  .rdata
			rid      => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rid,       --                  .rid
			rlast    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rlast,     --                  .rlast
			rready   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rready,    --                  .rready
			rresp    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rresp,     --                  .rresp
			rvalid   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rvalid,    --                  .rvalid
			wdata    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_wdata,     --                  .wdata
			wlast    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_wlast,     --                  .wlast
			wready   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_wready,    --                  .wready
			wstrb    => mm_interconnect_0_axi4slave_0_altera_axi4_slave_wstrb,     --                  .wstrb
			wvalid   => mm_interconnect_0_axi4slave_0_altera_axi4_slave_wvalid,    --                  .wvalid
			RST_N    => rst_controller_reset_out_reset_ports_inv                   --        reset_sink.reset_n
		);

	aximaster_0 : component Example3_axiMaster_0
		port map (
			CLK      => clk_clk,                                  --              clock.clk
			araddr   => aximaster_0_altera_axi4_master_araddr,    -- altera_axi4_master.araddr
			arburst  => aximaster_0_altera_axi4_master_arburst,   --                   .arburst
			arcache  => aximaster_0_altera_axi4_master_arcache,   --                   .arcache
			arid     => aximaster_0_altera_axi4_master_arid,      --                   .arid
			arlen    => aximaster_0_altera_axi4_master_arlen,     --                   .arlen
			arlock   => aximaster_0_altera_axi4_master_arlock,    --                   .arlock
			arprot   => aximaster_0_altera_axi4_master_arprot,    --                   .arprot
			arqos    => aximaster_0_altera_axi4_master_arqos,     --                   .arqos
			arready  => aximaster_0_altera_axi4_master_arready,   --                   .arready
			arregion => aximaster_0_altera_axi4_master_arregion,  --                   .arregion
			arsize   => aximaster_0_altera_axi4_master_arsize,    --                   .arsize
			arvalid  => aximaster_0_altera_axi4_master_arvalid,   --                   .arvalid
			awaddr   => aximaster_0_altera_axi4_master_awaddr,    --                   .awaddr
			awburst  => aximaster_0_altera_axi4_master_awburst,   --                   .awburst
			awcache  => aximaster_0_altera_axi4_master_awcache,   --                   .awcache
			awid     => aximaster_0_altera_axi4_master_awid,      --                   .awid
			awlen    => aximaster_0_altera_axi4_master_awlen,     --                   .awlen
			awlock   => aximaster_0_altera_axi4_master_awlock,    --                   .awlock
			awprot   => aximaster_0_altera_axi4_master_awprot,    --                   .awprot
			awqos    => aximaster_0_altera_axi4_master_awqos,     --                   .awqos
			awready  => aximaster_0_altera_axi4_master_awready,   --                   .awready
			awregion => aximaster_0_altera_axi4_master_awregion,  --                   .awregion
			awsize   => aximaster_0_altera_axi4_master_awsize,    --                   .awsize
			awvalid  => aximaster_0_altera_axi4_master_awvalid,   --                   .awvalid
			bid      => aximaster_0_altera_axi4_master_bid,       --                   .bid
			bready   => aximaster_0_altera_axi4_master_bready,    --                   .bready
			bresp    => aximaster_0_altera_axi4_master_bresp,     --                   .bresp
			bvalid   => aximaster_0_altera_axi4_master_bvalid,    --                   .bvalid
			rdata    => aximaster_0_altera_axi4_master_rdata,     --                   .rdata
			rid      => aximaster_0_altera_axi4_master_rid,       --                   .rid
			rlast    => aximaster_0_altera_axi4_master_rlast,     --                   .rlast
			rready   => aximaster_0_altera_axi4_master_rready,    --                   .rready
			rresp    => aximaster_0_altera_axi4_master_rresp,     --                   .rresp
			rvalid   => aximaster_0_altera_axi4_master_rvalid,    --                   .rvalid
			wdata    => aximaster_0_altera_axi4_master_wdata,     --                   .wdata
			wlast    => aximaster_0_altera_axi4_master_wlast,     --                   .wlast
			wready   => aximaster_0_altera_axi4_master_wready,    --                   .wready
			wstrb    => aximaster_0_altera_axi4_master_wstrb,     --                   .wstrb
			wvalid   => aximaster_0_altera_axi4_master_wvalid,    --                   .wvalid
			RST_N    => rst_controller_reset_out_reset_ports_inv  --         reset_sink.reset_n
		);

	mm_interconnect_0 : component Example3_mm_interconnect_0
		port map (
			axi4Slave_0_altera_axi4_slave_awid                 => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awid,     --                axi4Slave_0_altera_axi4_slave.awid
			axi4Slave_0_altera_axi4_slave_awaddr               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awaddr,   --                                             .awaddr
			axi4Slave_0_altera_axi4_slave_awlen                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awlen,    --                                             .awlen
			axi4Slave_0_altera_axi4_slave_awsize               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awsize,   --                                             .awsize
			axi4Slave_0_altera_axi4_slave_awburst              => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awburst,  --                                             .awburst
			axi4Slave_0_altera_axi4_slave_awlock               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awlock,   --                                             .awlock
			axi4Slave_0_altera_axi4_slave_awcache              => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awcache,  --                                             .awcache
			axi4Slave_0_altera_axi4_slave_awprot               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awprot,   --                                             .awprot
			axi4Slave_0_altera_axi4_slave_awqos                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awqos,    --                                             .awqos
			axi4Slave_0_altera_axi4_slave_awregion             => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awregion, --                                             .awregion
			axi4Slave_0_altera_axi4_slave_awvalid              => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awvalid,  --                                             .awvalid
			axi4Slave_0_altera_axi4_slave_awready              => mm_interconnect_0_axi4slave_0_altera_axi4_slave_awready,  --                                             .awready
			axi4Slave_0_altera_axi4_slave_wdata                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_wdata,    --                                             .wdata
			axi4Slave_0_altera_axi4_slave_wstrb                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_wstrb,    --                                             .wstrb
			axi4Slave_0_altera_axi4_slave_wlast                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_wlast,    --                                             .wlast
			axi4Slave_0_altera_axi4_slave_wvalid               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_wvalid,   --                                             .wvalid
			axi4Slave_0_altera_axi4_slave_wready               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_wready,   --                                             .wready
			axi4Slave_0_altera_axi4_slave_bid                  => mm_interconnect_0_axi4slave_0_altera_axi4_slave_bid,      --                                             .bid
			axi4Slave_0_altera_axi4_slave_bresp                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_bresp,    --                                             .bresp
			axi4Slave_0_altera_axi4_slave_bvalid               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_bvalid,   --                                             .bvalid
			axi4Slave_0_altera_axi4_slave_bready               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_bready,   --                                             .bready
			axi4Slave_0_altera_axi4_slave_arid                 => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arid,     --                                             .arid
			axi4Slave_0_altera_axi4_slave_araddr               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_araddr,   --                                             .araddr
			axi4Slave_0_altera_axi4_slave_arlen                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arlen,    --                                             .arlen
			axi4Slave_0_altera_axi4_slave_arsize               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arsize,   --                                             .arsize
			axi4Slave_0_altera_axi4_slave_arburst              => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arburst,  --                                             .arburst
			axi4Slave_0_altera_axi4_slave_arlock               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arlock,   --                                             .arlock
			axi4Slave_0_altera_axi4_slave_arcache              => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arcache,  --                                             .arcache
			axi4Slave_0_altera_axi4_slave_arprot               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arprot,   --                                             .arprot
			axi4Slave_0_altera_axi4_slave_arqos                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arqos,    --                                             .arqos
			axi4Slave_0_altera_axi4_slave_arregion             => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arregion, --                                             .arregion
			axi4Slave_0_altera_axi4_slave_arvalid              => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arvalid,  --                                             .arvalid
			axi4Slave_0_altera_axi4_slave_arready              => mm_interconnect_0_axi4slave_0_altera_axi4_slave_arready,  --                                             .arready
			axi4Slave_0_altera_axi4_slave_rid                  => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rid,      --                                             .rid
			axi4Slave_0_altera_axi4_slave_rdata                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rdata,    --                                             .rdata
			axi4Slave_0_altera_axi4_slave_rresp                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rresp,    --                                             .rresp
			axi4Slave_0_altera_axi4_slave_rlast                => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rlast,    --                                             .rlast
			axi4Slave_0_altera_axi4_slave_rvalid               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rvalid,   --                                             .rvalid
			axi4Slave_0_altera_axi4_slave_rready               => mm_interconnect_0_axi4slave_0_altera_axi4_slave_rready,   --                                             .rready
			axiMaster_0_altera_axi4_master_awid(0)             => aximaster_0_altera_axi4_master_awid,                      --               axiMaster_0_altera_axi4_master.awid
			axiMaster_0_altera_axi4_master_awaddr              => aximaster_0_altera_axi4_master_awaddr,                    --                                             .awaddr
			axiMaster_0_altera_axi4_master_awlen               => aximaster_0_altera_axi4_master_awlen,                     --                                             .awlen
			axiMaster_0_altera_axi4_master_awsize              => aximaster_0_altera_axi4_master_awsize,                    --                                             .awsize
			axiMaster_0_altera_axi4_master_awburst             => aximaster_0_altera_axi4_master_awburst,                   --                                             .awburst
			axiMaster_0_altera_axi4_master_awlock(0)           => aximaster_0_altera_axi4_master_awlock,                    --                                             .awlock
			axiMaster_0_altera_axi4_master_awcache             => aximaster_0_altera_axi4_master_awcache,                   --                                             .awcache
			axiMaster_0_altera_axi4_master_awprot              => aximaster_0_altera_axi4_master_awprot,                    --                                             .awprot
			axiMaster_0_altera_axi4_master_awqos               => aximaster_0_altera_axi4_master_awqos,                     --                                             .awqos
			axiMaster_0_altera_axi4_master_awregion            => aximaster_0_altera_axi4_master_awregion,                  --                                             .awregion
			axiMaster_0_altera_axi4_master_awvalid             => aximaster_0_altera_axi4_master_awvalid,                   --                                             .awvalid
			axiMaster_0_altera_axi4_master_awready             => aximaster_0_altera_axi4_master_awready,                   --                                             .awready
			axiMaster_0_altera_axi4_master_wdata               => aximaster_0_altera_axi4_master_wdata,                     --                                             .wdata
			axiMaster_0_altera_axi4_master_wstrb               => aximaster_0_altera_axi4_master_wstrb,                     --                                             .wstrb
			axiMaster_0_altera_axi4_master_wlast               => aximaster_0_altera_axi4_master_wlast,                     --                                             .wlast
			axiMaster_0_altera_axi4_master_wvalid              => aximaster_0_altera_axi4_master_wvalid,                    --                                             .wvalid
			axiMaster_0_altera_axi4_master_wready              => aximaster_0_altera_axi4_master_wready,                    --                                             .wready
			axiMaster_0_altera_axi4_master_bid(0)              => aximaster_0_altera_axi4_master_bid,                       --                                             .bid
			axiMaster_0_altera_axi4_master_bresp               => aximaster_0_altera_axi4_master_bresp,                     --                                             .bresp
			axiMaster_0_altera_axi4_master_bvalid              => aximaster_0_altera_axi4_master_bvalid,                    --                                             .bvalid
			axiMaster_0_altera_axi4_master_bready              => aximaster_0_altera_axi4_master_bready,                    --                                             .bready
			axiMaster_0_altera_axi4_master_arid(0)             => aximaster_0_altera_axi4_master_arid,                      --                                             .arid
			axiMaster_0_altera_axi4_master_araddr              => aximaster_0_altera_axi4_master_araddr,                    --                                             .araddr
			axiMaster_0_altera_axi4_master_arlen               => aximaster_0_altera_axi4_master_arlen,                     --                                             .arlen
			axiMaster_0_altera_axi4_master_arsize              => aximaster_0_altera_axi4_master_arsize,                    --                                             .arsize
			axiMaster_0_altera_axi4_master_arburst             => aximaster_0_altera_axi4_master_arburst,                   --                                             .arburst
			axiMaster_0_altera_axi4_master_arlock(0)           => aximaster_0_altera_axi4_master_arlock,                    --                                             .arlock
			axiMaster_0_altera_axi4_master_arcache             => aximaster_0_altera_axi4_master_arcache,                   --                                             .arcache
			axiMaster_0_altera_axi4_master_arprot              => aximaster_0_altera_axi4_master_arprot,                    --                                             .arprot
			axiMaster_0_altera_axi4_master_arqos               => aximaster_0_altera_axi4_master_arqos,                     --                                             .arqos
			axiMaster_0_altera_axi4_master_arregion            => aximaster_0_altera_axi4_master_arregion,                  --                                             .arregion
			axiMaster_0_altera_axi4_master_arvalid             => aximaster_0_altera_axi4_master_arvalid,                   --                                             .arvalid
			axiMaster_0_altera_axi4_master_arready             => aximaster_0_altera_axi4_master_arready,                   --                                             .arready
			axiMaster_0_altera_axi4_master_rid(0)              => aximaster_0_altera_axi4_master_rid,                       --                                             .rid
			axiMaster_0_altera_axi4_master_rdata               => aximaster_0_altera_axi4_master_rdata,                     --                                             .rdata
			axiMaster_0_altera_axi4_master_rresp               => aximaster_0_altera_axi4_master_rresp,                     --                                             .rresp
			axiMaster_0_altera_axi4_master_rlast               => aximaster_0_altera_axi4_master_rlast,                     --                                             .rlast
			axiMaster_0_altera_axi4_master_rvalid              => aximaster_0_altera_axi4_master_rvalid,                    --                                             .rvalid
			axiMaster_0_altera_axi4_master_rready              => aximaster_0_altera_axi4_master_rready,                    --                                             .rready
			clk_0_clk_clk                                      => clk_clk,                                                  --                                    clk_0_clk.clk
			axiMaster_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset                            -- axiMaster_0_reset_sink_reset_bridge_in_reset.reset
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of Example3
