// Example3.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module Example3 (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire    [1:0] axi4master2_0_altera_axi4_master_awburst;                  // axi4Master2_0:awburst -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awburst
	wire    [3:0] axi4master2_0_altera_axi4_master_arregion;                 // axi4Master2_0:arregion -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_arregion
	wire    [7:0] axi4master2_0_altera_axi4_master_arlen;                    // axi4Master2_0:arlen -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_arlen
	wire    [3:0] axi4master2_0_altera_axi4_master_arqos;                    // axi4Master2_0:arqos -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_arqos
	wire          axi4master2_0_altera_axi4_master_wready;                   // mm_interconnect_0:axi4Master2_0_altera_axi4_master_wready -> axi4Master2_0:wready
	wire   [15:0] axi4master2_0_altera_axi4_master_wstrb;                    // axi4Master2_0:wstrb -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_wstrb
	wire          axi4master2_0_altera_axi4_master_rid;                      // mm_interconnect_0:axi4Master2_0_altera_axi4_master_rid -> axi4Master2_0:rid
	wire          axi4master2_0_altera_axi4_master_rready;                   // axi4Master2_0:rready -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_rready
	wire    [7:0] axi4master2_0_altera_axi4_master_awlen;                    // axi4Master2_0:awlen -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awlen
	wire    [3:0] axi4master2_0_altera_axi4_master_awqos;                    // axi4Master2_0:awqos -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awqos
	wire    [3:0] axi4master2_0_altera_axi4_master_arcache;                  // axi4Master2_0:arcache -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_arcache
	wire   [13:0] axi4master2_0_altera_axi4_master_araddr;                   // axi4Master2_0:araddr -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_araddr
	wire          axi4master2_0_altera_axi4_master_wvalid;                   // axi4Master2_0:wvalid -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_wvalid
	wire    [2:0] axi4master2_0_altera_axi4_master_arprot;                   // axi4Master2_0:arprot -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_arprot
	wire          axi4master2_0_altera_axi4_master_arvalid;                  // axi4Master2_0:arvalid -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_arvalid
	wire    [2:0] axi4master2_0_altera_axi4_master_awprot;                   // axi4Master2_0:awprot -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awprot
	wire  [127:0] axi4master2_0_altera_axi4_master_wdata;                    // axi4Master2_0:wdata -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_wdata
	wire          axi4master2_0_altera_axi4_master_arid;                     // axi4Master2_0:arid -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_arid
	wire    [3:0] axi4master2_0_altera_axi4_master_awcache;                  // axi4Master2_0:awcache -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awcache
	wire          axi4master2_0_altera_axi4_master_arlock;                   // axi4Master2_0:arlock -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_arlock
	wire          axi4master2_0_altera_axi4_master_awlock;                   // axi4Master2_0:awlock -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awlock
	wire   [13:0] axi4master2_0_altera_axi4_master_awaddr;                   // axi4Master2_0:awaddr -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awaddr
	wire          axi4master2_0_altera_axi4_master_arready;                  // mm_interconnect_0:axi4Master2_0_altera_axi4_master_arready -> axi4Master2_0:arready
	wire    [1:0] axi4master2_0_altera_axi4_master_bresp;                    // mm_interconnect_0:axi4Master2_0_altera_axi4_master_bresp -> axi4Master2_0:bresp
	wire  [127:0] axi4master2_0_altera_axi4_master_rdata;                    // mm_interconnect_0:axi4Master2_0_altera_axi4_master_rdata -> axi4Master2_0:rdata
	wire    [1:0] axi4master2_0_altera_axi4_master_arburst;                  // axi4Master2_0:arburst -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_arburst
	wire          axi4master2_0_altera_axi4_master_awready;                  // mm_interconnect_0:axi4Master2_0_altera_axi4_master_awready -> axi4Master2_0:awready
	wire    [2:0] axi4master2_0_altera_axi4_master_arsize;                   // axi4Master2_0:arsize -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_arsize
	wire          axi4master2_0_altera_axi4_master_bready;                   // axi4Master2_0:bready -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_bready
	wire          axi4master2_0_altera_axi4_master_rlast;                    // mm_interconnect_0:axi4Master2_0_altera_axi4_master_rlast -> axi4Master2_0:rlast
	wire          axi4master2_0_altera_axi4_master_wlast;                    // axi4Master2_0:wlast -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_wlast
	wire    [3:0] axi4master2_0_altera_axi4_master_awregion;                 // axi4Master2_0:awregion -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awregion
	wire    [1:0] axi4master2_0_altera_axi4_master_rresp;                    // mm_interconnect_0:axi4Master2_0_altera_axi4_master_rresp -> axi4Master2_0:rresp
	wire          axi4master2_0_altera_axi4_master_awid;                     // axi4Master2_0:awid -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awid
	wire          axi4master2_0_altera_axi4_master_bid;                      // mm_interconnect_0:axi4Master2_0_altera_axi4_master_bid -> axi4Master2_0:bid
	wire          axi4master2_0_altera_axi4_master_bvalid;                   // mm_interconnect_0:axi4Master2_0_altera_axi4_master_bvalid -> axi4Master2_0:bvalid
	wire    [2:0] axi4master2_0_altera_axi4_master_awsize;                   // axi4Master2_0:awsize -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awsize
	wire          axi4master2_0_altera_axi4_master_awvalid;                  // axi4Master2_0:awvalid -> mm_interconnect_0:axi4Master2_0_altera_axi4_master_awvalid
	wire          axi4master2_0_altera_axi4_master_rvalid;                   // mm_interconnect_0:axi4Master2_0_altera_axi4_master_rvalid -> axi4Master2_0:rvalid
	wire    [1:0] axi4master1_0_altera_axi4_master_awburst;                  // axi4Master1_0:awburst -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awburst
	wire    [3:0] axi4master1_0_altera_axi4_master_arregion;                 // axi4Master1_0:arregion -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_arregion
	wire    [7:0] axi4master1_0_altera_axi4_master_arlen;                    // axi4Master1_0:arlen -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_arlen
	wire    [3:0] axi4master1_0_altera_axi4_master_arqos;                    // axi4Master1_0:arqos -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_arqos
	wire          axi4master1_0_altera_axi4_master_wready;                   // mm_interconnect_0:axi4Master1_0_altera_axi4_master_wready -> axi4Master1_0:wready
	wire   [15:0] axi4master1_0_altera_axi4_master_wstrb;                    // axi4Master1_0:wstrb -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_wstrb
	wire          axi4master1_0_altera_axi4_master_rid;                      // mm_interconnect_0:axi4Master1_0_altera_axi4_master_rid -> axi4Master1_0:rid
	wire          axi4master1_0_altera_axi4_master_rready;                   // axi4Master1_0:rready -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_rready
	wire    [7:0] axi4master1_0_altera_axi4_master_awlen;                    // axi4Master1_0:awlen -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awlen
	wire    [3:0] axi4master1_0_altera_axi4_master_awqos;                    // axi4Master1_0:awqos -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awqos
	wire    [3:0] axi4master1_0_altera_axi4_master_arcache;                  // axi4Master1_0:arcache -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_arcache
	wire   [13:0] axi4master1_0_altera_axi4_master_araddr;                   // axi4Master1_0:araddr -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_araddr
	wire          axi4master1_0_altera_axi4_master_wvalid;                   // axi4Master1_0:wvalid -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_wvalid
	wire    [2:0] axi4master1_0_altera_axi4_master_arprot;                   // axi4Master1_0:arprot -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_arprot
	wire          axi4master1_0_altera_axi4_master_arvalid;                  // axi4Master1_0:arvalid -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_arvalid
	wire    [2:0] axi4master1_0_altera_axi4_master_awprot;                   // axi4Master1_0:awprot -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awprot
	wire  [127:0] axi4master1_0_altera_axi4_master_wdata;                    // axi4Master1_0:wdata -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_wdata
	wire          axi4master1_0_altera_axi4_master_arid;                     // axi4Master1_0:arid -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_arid
	wire    [3:0] axi4master1_0_altera_axi4_master_awcache;                  // axi4Master1_0:awcache -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awcache
	wire          axi4master1_0_altera_axi4_master_arlock;                   // axi4Master1_0:arlock -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_arlock
	wire          axi4master1_0_altera_axi4_master_awlock;                   // axi4Master1_0:awlock -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awlock
	wire   [13:0] axi4master1_0_altera_axi4_master_awaddr;                   // axi4Master1_0:awaddr -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awaddr
	wire          axi4master1_0_altera_axi4_master_arready;                  // mm_interconnect_0:axi4Master1_0_altera_axi4_master_arready -> axi4Master1_0:arready
	wire    [1:0] axi4master1_0_altera_axi4_master_bresp;                    // mm_interconnect_0:axi4Master1_0_altera_axi4_master_bresp -> axi4Master1_0:bresp
	wire  [127:0] axi4master1_0_altera_axi4_master_rdata;                    // mm_interconnect_0:axi4Master1_0_altera_axi4_master_rdata -> axi4Master1_0:rdata
	wire    [1:0] axi4master1_0_altera_axi4_master_arburst;                  // axi4Master1_0:arburst -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_arburst
	wire          axi4master1_0_altera_axi4_master_awready;                  // mm_interconnect_0:axi4Master1_0_altera_axi4_master_awready -> axi4Master1_0:awready
	wire    [2:0] axi4master1_0_altera_axi4_master_arsize;                   // axi4Master1_0:arsize -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_arsize
	wire          axi4master1_0_altera_axi4_master_bready;                   // axi4Master1_0:bready -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_bready
	wire          axi4master1_0_altera_axi4_master_rlast;                    // mm_interconnect_0:axi4Master1_0_altera_axi4_master_rlast -> axi4Master1_0:rlast
	wire          axi4master1_0_altera_axi4_master_wlast;                    // axi4Master1_0:wlast -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_wlast
	wire    [3:0] axi4master1_0_altera_axi4_master_awregion;                 // axi4Master1_0:awregion -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awregion
	wire    [1:0] axi4master1_0_altera_axi4_master_rresp;                    // mm_interconnect_0:axi4Master1_0_altera_axi4_master_rresp -> axi4Master1_0:rresp
	wire          axi4master1_0_altera_axi4_master_awid;                     // axi4Master1_0:awid -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awid
	wire          axi4master1_0_altera_axi4_master_bid;                      // mm_interconnect_0:axi4Master1_0_altera_axi4_master_bid -> axi4Master1_0:bid
	wire          axi4master1_0_altera_axi4_master_bvalid;                   // mm_interconnect_0:axi4Master1_0_altera_axi4_master_bvalid -> axi4Master1_0:bvalid
	wire    [2:0] axi4master1_0_altera_axi4_master_awsize;                   // axi4Master1_0:awsize -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awsize
	wire          axi4master1_0_altera_axi4_master_awvalid;                  // axi4Master1_0:awvalid -> mm_interconnect_0:axi4Master1_0_altera_axi4_master_awvalid
	wire          axi4master1_0_altera_axi4_master_rvalid;                   // mm_interconnect_0:axi4Master1_0_altera_axi4_master_rvalid -> axi4Master1_0:rvalid
	wire    [1:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awburst;  // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awburst -> axi4Slave5_0:awburst
	wire    [3:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arregion; // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arregion -> axi4Slave5_0:arregion
	wire    [7:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arlen;    // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arlen -> axi4Slave5_0:arlen
	wire    [3:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arqos;    // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arqos -> axi4Slave5_0:arqos
	wire   [15:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wstrb;    // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_wstrb -> axi4Slave5_0:wstrb
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wready;   // axi4Slave5_0:wready -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_wready
	wire    [1:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rid;      // axi4Slave5_0:rid -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_rid
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rready;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_rready -> axi4Slave5_0:rready
	wire    [7:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awlen;    // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awlen -> axi4Slave5_0:awlen
	wire    [3:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awqos;    // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awqos -> axi4Slave5_0:awqos
	wire    [3:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arcache;  // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arcache -> axi4Slave5_0:arcache
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wvalid;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_wvalid -> axi4Slave5_0:wvalid
	wire   [12:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_araddr;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_araddr -> axi4Slave5_0:araddr
	wire    [2:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arprot;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arprot -> axi4Slave5_0:arprot
	wire    [2:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awprot;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awprot -> axi4Slave5_0:awprot
	wire  [127:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wdata;    // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_wdata -> axi4Slave5_0:wdata
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arvalid;  // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arvalid -> axi4Slave5_0:arvalid
	wire    [3:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awcache;  // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awcache -> axi4Slave5_0:awcache
	wire    [1:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arid;     // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arid -> axi4Slave5_0:arid
	wire    [0:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arlock;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arlock -> axi4Slave5_0:arlock
	wire    [0:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awlock;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awlock -> axi4Slave5_0:awlock
	wire   [12:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awaddr;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awaddr -> axi4Slave5_0:awaddr
	wire    [1:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bresp;    // axi4Slave5_0:bresp -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_bresp
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arready;  // axi4Slave5_0:arready -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arready
	wire  [127:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rdata;    // axi4Slave5_0:rdata -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_rdata
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awready;  // axi4Slave5_0:awready -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awready
	wire    [1:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arburst;  // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arburst -> axi4Slave5_0:arburst
	wire    [2:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arsize;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_arsize -> axi4Slave5_0:arsize
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bready;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_bready -> axi4Slave5_0:bready
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rlast;    // axi4Slave5_0:rlast -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_rlast
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wlast;    // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_wlast -> axi4Slave5_0:wlast
	wire    [3:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awregion; // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awregion -> axi4Slave5_0:awregion
	wire    [1:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rresp;    // axi4Slave5_0:rresp -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_rresp
	wire    [1:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awid;     // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awid -> axi4Slave5_0:awid
	wire    [1:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bid;      // axi4Slave5_0:bid -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_bid
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bvalid;   // axi4Slave5_0:bvalid -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_bvalid
	wire    [2:0] mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awsize;   // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awsize -> axi4Slave5_0:awsize
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awvalid;  // mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_awvalid -> axi4Slave5_0:awvalid
	wire          mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rvalid;   // axi4Slave5_0:rvalid -> mm_interconnect_0:axi4Slave5_0_altera_axi4_slave_rvalid
	wire    [1:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awburst;  // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awburst -> axi4Slave7_0:awburst
	wire    [3:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arregion; // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arregion -> axi4Slave7_0:arregion
	wire    [7:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arlen;    // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arlen -> axi4Slave7_0:arlen
	wire    [3:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arqos;    // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arqos -> axi4Slave7_0:arqos
	wire   [15:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wstrb;    // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_wstrb -> axi4Slave7_0:wstrb
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wready;   // axi4Slave7_0:wready -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_wready
	wire    [1:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rid;      // axi4Slave7_0:rid -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_rid
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rready;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_rready -> axi4Slave7_0:rready
	wire    [7:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awlen;    // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awlen -> axi4Slave7_0:awlen
	wire    [3:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awqos;    // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awqos -> axi4Slave7_0:awqos
	wire    [3:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arcache;  // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arcache -> axi4Slave7_0:arcache
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wvalid;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_wvalid -> axi4Slave7_0:wvalid
	wire   [12:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_araddr;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_araddr -> axi4Slave7_0:araddr
	wire    [2:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arprot;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arprot -> axi4Slave7_0:arprot
	wire    [2:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awprot;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awprot -> axi4Slave7_0:awprot
	wire  [127:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wdata;    // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_wdata -> axi4Slave7_0:wdata
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arvalid;  // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arvalid -> axi4Slave7_0:arvalid
	wire    [3:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awcache;  // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awcache -> axi4Slave7_0:awcache
	wire    [1:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arid;     // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arid -> axi4Slave7_0:arid
	wire    [0:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arlock;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arlock -> axi4Slave7_0:arlock
	wire    [0:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awlock;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awlock -> axi4Slave7_0:awlock
	wire   [12:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awaddr;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awaddr -> axi4Slave7_0:awaddr
	wire    [1:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bresp;    // axi4Slave7_0:bresp -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_bresp
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arready;  // axi4Slave7_0:arready -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arready
	wire  [127:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rdata;    // axi4Slave7_0:rdata -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_rdata
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awready;  // axi4Slave7_0:awready -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awready
	wire    [1:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arburst;  // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arburst -> axi4Slave7_0:arburst
	wire    [2:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arsize;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_arsize -> axi4Slave7_0:arsize
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bready;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_bready -> axi4Slave7_0:bready
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rlast;    // axi4Slave7_0:rlast -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_rlast
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wlast;    // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_wlast -> axi4Slave7_0:wlast
	wire    [3:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awregion; // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awregion -> axi4Slave7_0:awregion
	wire    [1:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rresp;    // axi4Slave7_0:rresp -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_rresp
	wire    [1:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awid;     // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awid -> axi4Slave7_0:awid
	wire    [1:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bid;      // axi4Slave7_0:bid -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_bid
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bvalid;   // axi4Slave7_0:bvalid -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_bvalid
	wire    [2:0] mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awsize;   // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awsize -> axi4Slave7_0:awsize
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awvalid;  // mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_awvalid -> axi4Slave7_0:awvalid
	wire          mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rvalid;   // axi4Slave7_0:rvalid -> mm_interconnect_0:axi4Slave7_0_altera_axi4_slave_rvalid
	wire          rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [axi4Master1_0:RST_N, axi4Master2_0:RST_N, axi4Slave5_0:RST_N, axi4Slave7_0:RST_N, mm_interconnect_0:axi4Master2_0_reset_sink_reset_bridge_in_reset_reset]

	axiMaster1_synth axi4master1_0 (
		.CLK      (clk_clk),                                   //              clock.clk
		.araddr   (axi4master1_0_altera_axi4_master_araddr),   // altera_axi4_master.araddr
		.arburst  (axi4master1_0_altera_axi4_master_arburst),  //                   .arburst
		.arcache  (axi4master1_0_altera_axi4_master_arcache),  //                   .arcache
		.arid     (axi4master1_0_altera_axi4_master_arid),     //                   .arid
		.arlen    (axi4master1_0_altera_axi4_master_arlen),    //                   .arlen
		.arlock   (axi4master1_0_altera_axi4_master_arlock),   //                   .arlock
		.arprot   (axi4master1_0_altera_axi4_master_arprot),   //                   .arprot
		.arqos    (axi4master1_0_altera_axi4_master_arqos),    //                   .arqos
		.arready  (axi4master1_0_altera_axi4_master_arready),  //                   .arready
		.arregion (axi4master1_0_altera_axi4_master_arregion), //                   .arregion
		.arsize   (axi4master1_0_altera_axi4_master_arsize),   //                   .arsize
		.arvalid  (axi4master1_0_altera_axi4_master_arvalid),  //                   .arvalid
		.awaddr   (axi4master1_0_altera_axi4_master_awaddr),   //                   .awaddr
		.awburst  (axi4master1_0_altera_axi4_master_awburst),  //                   .awburst
		.awcache  (axi4master1_0_altera_axi4_master_awcache),  //                   .awcache
		.awid     (axi4master1_0_altera_axi4_master_awid),     //                   .awid
		.awlen    (axi4master1_0_altera_axi4_master_awlen),    //                   .awlen
		.awlock   (axi4master1_0_altera_axi4_master_awlock),   //                   .awlock
		.awprot   (axi4master1_0_altera_axi4_master_awprot),   //                   .awprot
		.awqos    (axi4master1_0_altera_axi4_master_awqos),    //                   .awqos
		.awready  (axi4master1_0_altera_axi4_master_awready),  //                   .awready
		.awregion (axi4master1_0_altera_axi4_master_awregion), //                   .awregion
		.awsize   (axi4master1_0_altera_axi4_master_awsize),   //                   .awsize
		.awvalid  (axi4master1_0_altera_axi4_master_awvalid),  //                   .awvalid
		.bid      (axi4master1_0_altera_axi4_master_bid),      //                   .bid
		.bready   (axi4master1_0_altera_axi4_master_bready),   //                   .bready
		.bresp    (axi4master1_0_altera_axi4_master_bresp),    //                   .bresp
		.bvalid   (axi4master1_0_altera_axi4_master_bvalid),   //                   .bvalid
		.rdata    (axi4master1_0_altera_axi4_master_rdata),    //                   .rdata
		.rid      (axi4master1_0_altera_axi4_master_rid),      //                   .rid
		.rlast    (axi4master1_0_altera_axi4_master_rlast),    //                   .rlast
		.rready   (axi4master1_0_altera_axi4_master_rready),   //                   .rready
		.rresp    (axi4master1_0_altera_axi4_master_rresp),    //                   .rresp
		.rvalid   (axi4master1_0_altera_axi4_master_rvalid),   //                   .rvalid
		.wdata    (axi4master1_0_altera_axi4_master_wdata),    //                   .wdata
		.wlast    (axi4master1_0_altera_axi4_master_wlast),    //                   .wlast
		.wready   (axi4master1_0_altera_axi4_master_wready),   //                   .wready
		.wstrb    (axi4master1_0_altera_axi4_master_wstrb),    //                   .wstrb
		.wvalid   (axi4master1_0_altera_axi4_master_wvalid),   //                   .wvalid
		.RST_N    (~rst_controller_reset_out_reset)            //         reset_sink.reset_n
	);

	axiMaster2_synth axi4master2_0 (
		.CLK      (clk_clk),                                   //              clock.clk
		.araddr   (axi4master2_0_altera_axi4_master_araddr),   // altera_axi4_master.araddr
		.arburst  (axi4master2_0_altera_axi4_master_arburst),  //                   .arburst
		.arcache  (axi4master2_0_altera_axi4_master_arcache),  //                   .arcache
		.arid     (axi4master2_0_altera_axi4_master_arid),     //                   .arid
		.arlen    (axi4master2_0_altera_axi4_master_arlen),    //                   .arlen
		.arlock   (axi4master2_0_altera_axi4_master_arlock),   //                   .arlock
		.arprot   (axi4master2_0_altera_axi4_master_arprot),   //                   .arprot
		.arqos    (axi4master2_0_altera_axi4_master_arqos),    //                   .arqos
		.arready  (axi4master2_0_altera_axi4_master_arready),  //                   .arready
		.arregion (axi4master2_0_altera_axi4_master_arregion), //                   .arregion
		.arsize   (axi4master2_0_altera_axi4_master_arsize),   //                   .arsize
		.arvalid  (axi4master2_0_altera_axi4_master_arvalid),  //                   .arvalid
		.awaddr   (axi4master2_0_altera_axi4_master_awaddr),   //                   .awaddr
		.awburst  (axi4master2_0_altera_axi4_master_awburst),  //                   .awburst
		.awcache  (axi4master2_0_altera_axi4_master_awcache),  //                   .awcache
		.awid     (axi4master2_0_altera_axi4_master_awid),     //                   .awid
		.awlen    (axi4master2_0_altera_axi4_master_awlen),    //                   .awlen
		.awlock   (axi4master2_0_altera_axi4_master_awlock),   //                   .awlock
		.awprot   (axi4master2_0_altera_axi4_master_awprot),   //                   .awprot
		.awqos    (axi4master2_0_altera_axi4_master_awqos),    //                   .awqos
		.awready  (axi4master2_0_altera_axi4_master_awready),  //                   .awready
		.awregion (axi4master2_0_altera_axi4_master_awregion), //                   .awregion
		.awsize   (axi4master2_0_altera_axi4_master_awsize),   //                   .awsize
		.awvalid  (axi4master2_0_altera_axi4_master_awvalid),  //                   .awvalid
		.bid      (axi4master2_0_altera_axi4_master_bid),      //                   .bid
		.bready   (axi4master2_0_altera_axi4_master_bready),   //                   .bready
		.bresp    (axi4master2_0_altera_axi4_master_bresp),    //                   .bresp
		.bvalid   (axi4master2_0_altera_axi4_master_bvalid),   //                   .bvalid
		.rdata    (axi4master2_0_altera_axi4_master_rdata),    //                   .rdata
		.rid      (axi4master2_0_altera_axi4_master_rid),      //                   .rid
		.rlast    (axi4master2_0_altera_axi4_master_rlast),    //                   .rlast
		.rready   (axi4master2_0_altera_axi4_master_rready),   //                   .rready
		.rresp    (axi4master2_0_altera_axi4_master_rresp),    //                   .rresp
		.rvalid   (axi4master2_0_altera_axi4_master_rvalid),   //                   .rvalid
		.wdata    (axi4master2_0_altera_axi4_master_wdata),    //                   .wdata
		.wlast    (axi4master2_0_altera_axi4_master_wlast),    //                   .wlast
		.wready   (axi4master2_0_altera_axi4_master_wready),   //                   .wready
		.wstrb    (axi4master2_0_altera_axi4_master_wstrb),    //                   .wstrb
		.wvalid   (axi4master2_0_altera_axi4_master_wvalid),   //                   .wvalid
		.RST_N    (~rst_controller_reset_out_reset)            //         reset_sink.reset_n
	);

	axiSlave5_synth axi4slave5_0 (
		.CLK      (clk_clk),                                                   //             clock.clk
		.araddr   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_araddr),   // altera_axi4_slave.araddr
		.arburst  (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arburst),  //                  .arburst
		.arcache  (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arcache),  //                  .arcache
		.arid     (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arid),     //                  .arid
		.arlen    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arlen),    //                  .arlen
		.arlock   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arlock),   //                  .arlock
		.arprot   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arprot),   //                  .arprot
		.arqos    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arqos),    //                  .arqos
		.arready  (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arready),  //                  .arready
		.arregion (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arregion), //                  .arregion
		.arsize   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arsize),   //                  .arsize
		.arvalid  (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arvalid),  //                  .arvalid
		.awaddr   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awaddr),   //                  .awaddr
		.awburst  (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awburst),  //                  .awburst
		.awcache  (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awcache),  //                  .awcache
		.awid     (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awid),     //                  .awid
		.awlen    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awlen),    //                  .awlen
		.awlock   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awlock),   //                  .awlock
		.awprot   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awprot),   //                  .awprot
		.awqos    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awqos),    //                  .awqos
		.awready  (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awready),  //                  .awready
		.awregion (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awregion), //                  .awregion
		.awsize   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awsize),   //                  .awsize
		.awvalid  (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awvalid),  //                  .awvalid
		.bid      (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bid),      //                  .bid
		.bready   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bready),   //                  .bready
		.bresp    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bresp),    //                  .bresp
		.bvalid   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bvalid),   //                  .bvalid
		.rdata    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rdata),    //                  .rdata
		.rid      (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rid),      //                  .rid
		.rlast    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rlast),    //                  .rlast
		.rready   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rready),   //                  .rready
		.rresp    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rresp),    //                  .rresp
		.rvalid   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rvalid),   //                  .rvalid
		.wdata    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wdata),    //                  .wdata
		.wlast    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wlast),    //                  .wlast
		.wready   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wready),   //                  .wready
		.wstrb    (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wstrb),    //                  .wstrb
		.wvalid   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wvalid),   //                  .wvalid
		.RST_N    (~rst_controller_reset_out_reset)                            //        reset_sink.reset_n
	);

	axiSlave7_synth axi4slave7_0 (
		.CLK      (clk_clk),                                                   //             clock.clk
		.araddr   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_araddr),   // altera_axi4_slave.araddr
		.arburst  (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arburst),  //                  .arburst
		.arcache  (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arcache),  //                  .arcache
		.arid     (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arid),     //                  .arid
		.arlen    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arlen),    //                  .arlen
		.arlock   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arlock),   //                  .arlock
		.arprot   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arprot),   //                  .arprot
		.arqos    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arqos),    //                  .arqos
		.arready  (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arready),  //                  .arready
		.arregion (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arregion), //                  .arregion
		.arsize   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arsize),   //                  .arsize
		.arvalid  (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arvalid),  //                  .arvalid
		.awaddr   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awaddr),   //                  .awaddr
		.awburst  (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awburst),  //                  .awburst
		.awcache  (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awcache),  //                  .awcache
		.awid     (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awid),     //                  .awid
		.awlen    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awlen),    //                  .awlen
		.awlock   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awlock),   //                  .awlock
		.awprot   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awprot),   //                  .awprot
		.awqos    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awqos),    //                  .awqos
		.awready  (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awready),  //                  .awready
		.awregion (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awregion), //                  .awregion
		.awsize   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awsize),   //                  .awsize
		.awvalid  (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awvalid),  //                  .awvalid
		.bid      (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bid),      //                  .bid
		.bready   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bready),   //                  .bready
		.bresp    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bresp),    //                  .bresp
		.bvalid   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bvalid),   //                  .bvalid
		.rdata    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rdata),    //                  .rdata
		.rid      (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rid),      //                  .rid
		.rlast    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rlast),    //                  .rlast
		.rready   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rready),   //                  .rready
		.rresp    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rresp),    //                  .rresp
		.rvalid   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rvalid),   //                  .rvalid
		.wdata    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wdata),    //                  .wdata
		.wlast    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wlast),    //                  .wlast
		.wready   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wready),   //                  .wready
		.wstrb    (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wstrb),    //                  .wstrb
		.wvalid   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wvalid),   //                  .wvalid
		.RST_N    (~rst_controller_reset_out_reset)                            //        reset_sink.reset_n
	);

	Example3_mm_interconnect_0 mm_interconnect_0 (
		.axi4Master1_0_altera_axi4_master_awid                (axi4master1_0_altera_axi4_master_awid),                     //               axi4Master1_0_altera_axi4_master.awid
		.axi4Master1_0_altera_axi4_master_awaddr              (axi4master1_0_altera_axi4_master_awaddr),                   //                                               .awaddr
		.axi4Master1_0_altera_axi4_master_awlen               (axi4master1_0_altera_axi4_master_awlen),                    //                                               .awlen
		.axi4Master1_0_altera_axi4_master_awsize              (axi4master1_0_altera_axi4_master_awsize),                   //                                               .awsize
		.axi4Master1_0_altera_axi4_master_awburst             (axi4master1_0_altera_axi4_master_awburst),                  //                                               .awburst
		.axi4Master1_0_altera_axi4_master_awlock              (axi4master1_0_altera_axi4_master_awlock),                   //                                               .awlock
		.axi4Master1_0_altera_axi4_master_awcache             (axi4master1_0_altera_axi4_master_awcache),                  //                                               .awcache
		.axi4Master1_0_altera_axi4_master_awprot              (axi4master1_0_altera_axi4_master_awprot),                   //                                               .awprot
		.axi4Master1_0_altera_axi4_master_awqos               (axi4master1_0_altera_axi4_master_awqos),                    //                                               .awqos
		.axi4Master1_0_altera_axi4_master_awregion            (axi4master1_0_altera_axi4_master_awregion),                 //                                               .awregion
		.axi4Master1_0_altera_axi4_master_awvalid             (axi4master1_0_altera_axi4_master_awvalid),                  //                                               .awvalid
		.axi4Master1_0_altera_axi4_master_awready             (axi4master1_0_altera_axi4_master_awready),                  //                                               .awready
		.axi4Master1_0_altera_axi4_master_wdata               (axi4master1_0_altera_axi4_master_wdata),                    //                                               .wdata
		.axi4Master1_0_altera_axi4_master_wstrb               (axi4master1_0_altera_axi4_master_wstrb),                    //                                               .wstrb
		.axi4Master1_0_altera_axi4_master_wlast               (axi4master1_0_altera_axi4_master_wlast),                    //                                               .wlast
		.axi4Master1_0_altera_axi4_master_wvalid              (axi4master1_0_altera_axi4_master_wvalid),                   //                                               .wvalid
		.axi4Master1_0_altera_axi4_master_wready              (axi4master1_0_altera_axi4_master_wready),                   //                                               .wready
		.axi4Master1_0_altera_axi4_master_bid                 (axi4master1_0_altera_axi4_master_bid),                      //                                               .bid
		.axi4Master1_0_altera_axi4_master_bresp               (axi4master1_0_altera_axi4_master_bresp),                    //                                               .bresp
		.axi4Master1_0_altera_axi4_master_bvalid              (axi4master1_0_altera_axi4_master_bvalid),                   //                                               .bvalid
		.axi4Master1_0_altera_axi4_master_bready              (axi4master1_0_altera_axi4_master_bready),                   //                                               .bready
		.axi4Master1_0_altera_axi4_master_arid                (axi4master1_0_altera_axi4_master_arid),                     //                                               .arid
		.axi4Master1_0_altera_axi4_master_araddr              (axi4master1_0_altera_axi4_master_araddr),                   //                                               .araddr
		.axi4Master1_0_altera_axi4_master_arlen               (axi4master1_0_altera_axi4_master_arlen),                    //                                               .arlen
		.axi4Master1_0_altera_axi4_master_arsize              (axi4master1_0_altera_axi4_master_arsize),                   //                                               .arsize
		.axi4Master1_0_altera_axi4_master_arburst             (axi4master1_0_altera_axi4_master_arburst),                  //                                               .arburst
		.axi4Master1_0_altera_axi4_master_arlock              (axi4master1_0_altera_axi4_master_arlock),                   //                                               .arlock
		.axi4Master1_0_altera_axi4_master_arcache             (axi4master1_0_altera_axi4_master_arcache),                  //                                               .arcache
		.axi4Master1_0_altera_axi4_master_arprot              (axi4master1_0_altera_axi4_master_arprot),                   //                                               .arprot
		.axi4Master1_0_altera_axi4_master_arqos               (axi4master1_0_altera_axi4_master_arqos),                    //                                               .arqos
		.axi4Master1_0_altera_axi4_master_arregion            (axi4master1_0_altera_axi4_master_arregion),                 //                                               .arregion
		.axi4Master1_0_altera_axi4_master_arvalid             (axi4master1_0_altera_axi4_master_arvalid),                  //                                               .arvalid
		.axi4Master1_0_altera_axi4_master_arready             (axi4master1_0_altera_axi4_master_arready),                  //                                               .arready
		.axi4Master1_0_altera_axi4_master_rid                 (axi4master1_0_altera_axi4_master_rid),                      //                                               .rid
		.axi4Master1_0_altera_axi4_master_rdata               (axi4master1_0_altera_axi4_master_rdata),                    //                                               .rdata
		.axi4Master1_0_altera_axi4_master_rresp               (axi4master1_0_altera_axi4_master_rresp),                    //                                               .rresp
		.axi4Master1_0_altera_axi4_master_rlast               (axi4master1_0_altera_axi4_master_rlast),                    //                                               .rlast
		.axi4Master1_0_altera_axi4_master_rvalid              (axi4master1_0_altera_axi4_master_rvalid),                   //                                               .rvalid
		.axi4Master1_0_altera_axi4_master_rready              (axi4master1_0_altera_axi4_master_rready),                   //                                               .rready
		.axi4Master2_0_altera_axi4_master_awid                (axi4master2_0_altera_axi4_master_awid),                     //               axi4Master2_0_altera_axi4_master.awid
		.axi4Master2_0_altera_axi4_master_awaddr              (axi4master2_0_altera_axi4_master_awaddr),                   //                                               .awaddr
		.axi4Master2_0_altera_axi4_master_awlen               (axi4master2_0_altera_axi4_master_awlen),                    //                                               .awlen
		.axi4Master2_0_altera_axi4_master_awsize              (axi4master2_0_altera_axi4_master_awsize),                   //                                               .awsize
		.axi4Master2_0_altera_axi4_master_awburst             (axi4master2_0_altera_axi4_master_awburst),                  //                                               .awburst
		.axi4Master2_0_altera_axi4_master_awlock              (axi4master2_0_altera_axi4_master_awlock),                   //                                               .awlock
		.axi4Master2_0_altera_axi4_master_awcache             (axi4master2_0_altera_axi4_master_awcache),                  //                                               .awcache
		.axi4Master2_0_altera_axi4_master_awprot              (axi4master2_0_altera_axi4_master_awprot),                   //                                               .awprot
		.axi4Master2_0_altera_axi4_master_awqos               (axi4master2_0_altera_axi4_master_awqos),                    //                                               .awqos
		.axi4Master2_0_altera_axi4_master_awregion            (axi4master2_0_altera_axi4_master_awregion),                 //                                               .awregion
		.axi4Master2_0_altera_axi4_master_awvalid             (axi4master2_0_altera_axi4_master_awvalid),                  //                                               .awvalid
		.axi4Master2_0_altera_axi4_master_awready             (axi4master2_0_altera_axi4_master_awready),                  //                                               .awready
		.axi4Master2_0_altera_axi4_master_wdata               (axi4master2_0_altera_axi4_master_wdata),                    //                                               .wdata
		.axi4Master2_0_altera_axi4_master_wstrb               (axi4master2_0_altera_axi4_master_wstrb),                    //                                               .wstrb
		.axi4Master2_0_altera_axi4_master_wlast               (axi4master2_0_altera_axi4_master_wlast),                    //                                               .wlast
		.axi4Master2_0_altera_axi4_master_wvalid              (axi4master2_0_altera_axi4_master_wvalid),                   //                                               .wvalid
		.axi4Master2_0_altera_axi4_master_wready              (axi4master2_0_altera_axi4_master_wready),                   //                                               .wready
		.axi4Master2_0_altera_axi4_master_bid                 (axi4master2_0_altera_axi4_master_bid),                      //                                               .bid
		.axi4Master2_0_altera_axi4_master_bresp               (axi4master2_0_altera_axi4_master_bresp),                    //                                               .bresp
		.axi4Master2_0_altera_axi4_master_bvalid              (axi4master2_0_altera_axi4_master_bvalid),                   //                                               .bvalid
		.axi4Master2_0_altera_axi4_master_bready              (axi4master2_0_altera_axi4_master_bready),                   //                                               .bready
		.axi4Master2_0_altera_axi4_master_arid                (axi4master2_0_altera_axi4_master_arid),                     //                                               .arid
		.axi4Master2_0_altera_axi4_master_araddr              (axi4master2_0_altera_axi4_master_araddr),                   //                                               .araddr
		.axi4Master2_0_altera_axi4_master_arlen               (axi4master2_0_altera_axi4_master_arlen),                    //                                               .arlen
		.axi4Master2_0_altera_axi4_master_arsize              (axi4master2_0_altera_axi4_master_arsize),                   //                                               .arsize
		.axi4Master2_0_altera_axi4_master_arburst             (axi4master2_0_altera_axi4_master_arburst),                  //                                               .arburst
		.axi4Master2_0_altera_axi4_master_arlock              (axi4master2_0_altera_axi4_master_arlock),                   //                                               .arlock
		.axi4Master2_0_altera_axi4_master_arcache             (axi4master2_0_altera_axi4_master_arcache),                  //                                               .arcache
		.axi4Master2_0_altera_axi4_master_arprot              (axi4master2_0_altera_axi4_master_arprot),                   //                                               .arprot
		.axi4Master2_0_altera_axi4_master_arqos               (axi4master2_0_altera_axi4_master_arqos),                    //                                               .arqos
		.axi4Master2_0_altera_axi4_master_arregion            (axi4master2_0_altera_axi4_master_arregion),                 //                                               .arregion
		.axi4Master2_0_altera_axi4_master_arvalid             (axi4master2_0_altera_axi4_master_arvalid),                  //                                               .arvalid
		.axi4Master2_0_altera_axi4_master_arready             (axi4master2_0_altera_axi4_master_arready),                  //                                               .arready
		.axi4Master2_0_altera_axi4_master_rid                 (axi4master2_0_altera_axi4_master_rid),                      //                                               .rid
		.axi4Master2_0_altera_axi4_master_rdata               (axi4master2_0_altera_axi4_master_rdata),                    //                                               .rdata
		.axi4Master2_0_altera_axi4_master_rresp               (axi4master2_0_altera_axi4_master_rresp),                    //                                               .rresp
		.axi4Master2_0_altera_axi4_master_rlast               (axi4master2_0_altera_axi4_master_rlast),                    //                                               .rlast
		.axi4Master2_0_altera_axi4_master_rvalid              (axi4master2_0_altera_axi4_master_rvalid),                   //                                               .rvalid
		.axi4Master2_0_altera_axi4_master_rready              (axi4master2_0_altera_axi4_master_rready),                   //                                               .rready
		.axi4Slave5_0_altera_axi4_slave_awid                  (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awid),     //                 axi4Slave5_0_altera_axi4_slave.awid
		.axi4Slave5_0_altera_axi4_slave_awaddr                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awaddr),   //                                               .awaddr
		.axi4Slave5_0_altera_axi4_slave_awlen                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awlen),    //                                               .awlen
		.axi4Slave5_0_altera_axi4_slave_awsize                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awsize),   //                                               .awsize
		.axi4Slave5_0_altera_axi4_slave_awburst               (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awburst),  //                                               .awburst
		.axi4Slave5_0_altera_axi4_slave_awlock                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awlock),   //                                               .awlock
		.axi4Slave5_0_altera_axi4_slave_awcache               (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awcache),  //                                               .awcache
		.axi4Slave5_0_altera_axi4_slave_awprot                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awprot),   //                                               .awprot
		.axi4Slave5_0_altera_axi4_slave_awqos                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awqos),    //                                               .awqos
		.axi4Slave5_0_altera_axi4_slave_awregion              (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awregion), //                                               .awregion
		.axi4Slave5_0_altera_axi4_slave_awvalid               (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awvalid),  //                                               .awvalid
		.axi4Slave5_0_altera_axi4_slave_awready               (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_awready),  //                                               .awready
		.axi4Slave5_0_altera_axi4_slave_wdata                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wdata),    //                                               .wdata
		.axi4Slave5_0_altera_axi4_slave_wstrb                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wstrb),    //                                               .wstrb
		.axi4Slave5_0_altera_axi4_slave_wlast                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wlast),    //                                               .wlast
		.axi4Slave5_0_altera_axi4_slave_wvalid                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wvalid),   //                                               .wvalid
		.axi4Slave5_0_altera_axi4_slave_wready                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_wready),   //                                               .wready
		.axi4Slave5_0_altera_axi4_slave_bid                   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bid),      //                                               .bid
		.axi4Slave5_0_altera_axi4_slave_bresp                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bresp),    //                                               .bresp
		.axi4Slave5_0_altera_axi4_slave_bvalid                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bvalid),   //                                               .bvalid
		.axi4Slave5_0_altera_axi4_slave_bready                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_bready),   //                                               .bready
		.axi4Slave5_0_altera_axi4_slave_arid                  (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arid),     //                                               .arid
		.axi4Slave5_0_altera_axi4_slave_araddr                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_araddr),   //                                               .araddr
		.axi4Slave5_0_altera_axi4_slave_arlen                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arlen),    //                                               .arlen
		.axi4Slave5_0_altera_axi4_slave_arsize                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arsize),   //                                               .arsize
		.axi4Slave5_0_altera_axi4_slave_arburst               (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arburst),  //                                               .arburst
		.axi4Slave5_0_altera_axi4_slave_arlock                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arlock),   //                                               .arlock
		.axi4Slave5_0_altera_axi4_slave_arcache               (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arcache),  //                                               .arcache
		.axi4Slave5_0_altera_axi4_slave_arprot                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arprot),   //                                               .arprot
		.axi4Slave5_0_altera_axi4_slave_arqos                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arqos),    //                                               .arqos
		.axi4Slave5_0_altera_axi4_slave_arregion              (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arregion), //                                               .arregion
		.axi4Slave5_0_altera_axi4_slave_arvalid               (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arvalid),  //                                               .arvalid
		.axi4Slave5_0_altera_axi4_slave_arready               (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_arready),  //                                               .arready
		.axi4Slave5_0_altera_axi4_slave_rid                   (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rid),      //                                               .rid
		.axi4Slave5_0_altera_axi4_slave_rdata                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rdata),    //                                               .rdata
		.axi4Slave5_0_altera_axi4_slave_rresp                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rresp),    //                                               .rresp
		.axi4Slave5_0_altera_axi4_slave_rlast                 (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rlast),    //                                               .rlast
		.axi4Slave5_0_altera_axi4_slave_rvalid                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rvalid),   //                                               .rvalid
		.axi4Slave5_0_altera_axi4_slave_rready                (mm_interconnect_0_axi4slave5_0_altera_axi4_slave_rready),   //                                               .rready
		.axi4Slave7_0_altera_axi4_slave_awid                  (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awid),     //                 axi4Slave7_0_altera_axi4_slave.awid
		.axi4Slave7_0_altera_axi4_slave_awaddr                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awaddr),   //                                               .awaddr
		.axi4Slave7_0_altera_axi4_slave_awlen                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awlen),    //                                               .awlen
		.axi4Slave7_0_altera_axi4_slave_awsize                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awsize),   //                                               .awsize
		.axi4Slave7_0_altera_axi4_slave_awburst               (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awburst),  //                                               .awburst
		.axi4Slave7_0_altera_axi4_slave_awlock                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awlock),   //                                               .awlock
		.axi4Slave7_0_altera_axi4_slave_awcache               (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awcache),  //                                               .awcache
		.axi4Slave7_0_altera_axi4_slave_awprot                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awprot),   //                                               .awprot
		.axi4Slave7_0_altera_axi4_slave_awqos                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awqos),    //                                               .awqos
		.axi4Slave7_0_altera_axi4_slave_awregion              (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awregion), //                                               .awregion
		.axi4Slave7_0_altera_axi4_slave_awvalid               (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awvalid),  //                                               .awvalid
		.axi4Slave7_0_altera_axi4_slave_awready               (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_awready),  //                                               .awready
		.axi4Slave7_0_altera_axi4_slave_wdata                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wdata),    //                                               .wdata
		.axi4Slave7_0_altera_axi4_slave_wstrb                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wstrb),    //                                               .wstrb
		.axi4Slave7_0_altera_axi4_slave_wlast                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wlast),    //                                               .wlast
		.axi4Slave7_0_altera_axi4_slave_wvalid                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wvalid),   //                                               .wvalid
		.axi4Slave7_0_altera_axi4_slave_wready                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_wready),   //                                               .wready
		.axi4Slave7_0_altera_axi4_slave_bid                   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bid),      //                                               .bid
		.axi4Slave7_0_altera_axi4_slave_bresp                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bresp),    //                                               .bresp
		.axi4Slave7_0_altera_axi4_slave_bvalid                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bvalid),   //                                               .bvalid
		.axi4Slave7_0_altera_axi4_slave_bready                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_bready),   //                                               .bready
		.axi4Slave7_0_altera_axi4_slave_arid                  (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arid),     //                                               .arid
		.axi4Slave7_0_altera_axi4_slave_araddr                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_araddr),   //                                               .araddr
		.axi4Slave7_0_altera_axi4_slave_arlen                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arlen),    //                                               .arlen
		.axi4Slave7_0_altera_axi4_slave_arsize                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arsize),   //                                               .arsize
		.axi4Slave7_0_altera_axi4_slave_arburst               (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arburst),  //                                               .arburst
		.axi4Slave7_0_altera_axi4_slave_arlock                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arlock),   //                                               .arlock
		.axi4Slave7_0_altera_axi4_slave_arcache               (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arcache),  //                                               .arcache
		.axi4Slave7_0_altera_axi4_slave_arprot                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arprot),   //                                               .arprot
		.axi4Slave7_0_altera_axi4_slave_arqos                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arqos),    //                                               .arqos
		.axi4Slave7_0_altera_axi4_slave_arregion              (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arregion), //                                               .arregion
		.axi4Slave7_0_altera_axi4_slave_arvalid               (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arvalid),  //                                               .arvalid
		.axi4Slave7_0_altera_axi4_slave_arready               (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_arready),  //                                               .arready
		.axi4Slave7_0_altera_axi4_slave_rid                   (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rid),      //                                               .rid
		.axi4Slave7_0_altera_axi4_slave_rdata                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rdata),    //                                               .rdata
		.axi4Slave7_0_altera_axi4_slave_rresp                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rresp),    //                                               .rresp
		.axi4Slave7_0_altera_axi4_slave_rlast                 (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rlast),    //                                               .rlast
		.axi4Slave7_0_altera_axi4_slave_rvalid                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rvalid),   //                                               .rvalid
		.axi4Slave7_0_altera_axi4_slave_rready                (mm_interconnect_0_axi4slave7_0_altera_axi4_slave_rready),   //                                               .rready
		.clk_0_clk_clk                                        (clk_clk),                                                   //                                      clk_0_clk.clk
		.axi4Master2_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset)                             // axi4Master2_0_reset_sink_reset_bridge_in_reset.reset
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
