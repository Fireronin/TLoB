package fifoChain;
// necessary packages
import GetPut::*;
import MemUtils::*;
import AXI4_Interconnect::*;
import FIFO::*;
import Core::*;
import Connectable::*;
// imported packages
import GPR_RegFile::*;
import AXI4_AR_Utils::*;
import CPU_Stage2::*;
import AXI4_Events_BitVectorable_Instance::*;
import DM_CPU_Req_Rsp::*;
import Prelude::*;
import AXI4_AXI4Lite_Bridges::*;
import AXI4::*;
import DM_Run_Control::*;
import PreludeBSV::*;
import Map::*;
import SpecialWires::*;
import MasterSlave::*;
import FF::*;
import CPU_Stage1::*;
import FixedPoint::*;
import RISCV_MBox::*;
import BUtils::*;
import Near_Mem_Caches::*;
import AXI::*;
import AXI4Lite_AR_Utils::*;
import GenerateHPMVector::*;
import AXI4Lite_AW_Utils::*;
import AXI4Stream_Types::*;
import Printf::*;
import DM_Abstract_Commands::*;
import Reserved::*;
import TLB::*;
import List::*;
import RegFile::*;
import ISA_Decls::*;
import ByteLane::*;
import Divide::*;
import SourceSink::*;
import CPU_StageD::*;
import Interconnect::*;
import DefaultValue::*;
import FIFOF_::*;
import Real::*;
import CacheCore::*;
import AXI4Lite::*;
import VnD::*;
import FPU::*;
import Debug::*;
import BlueUtils::*;
import AXI_Helpers::*;
import Array::*;
import RevertingVirtualReg::*;
import BuildVector::*;
import ToString::*;
import FIFOF::*;
import Vector::*;
import AXI4_W_Utils::*;
import CPU::*;
import TV_Taps::*;
import Memory::*;
import MemTypes::*;
import FBox_Top::*;
import UGFFFullOfUniqueInts::*;
import FIFOLevel::*;
import CSR_MIP::*;
import RoutableCHERI::*;
import AXI4_R_Utils::*;
import TurboFIFO::*;
import TwoWayBus::*;
import CSR_MSTATUS::*;
import TV_Info::*;
import Inout::*;
import SoC_Map::*;
import AXI4Lite_Interconnect::*;
import StatCounters::*;
import PLIC_16_2_7::*;
import ConfigReg::*;
import Branch_Predictor::*;
import CPU_Stage3::*;
import PerformanceMonitor::*;
import AXI4_Utils::*;
import EX_ALU_functions::*;
import SimpleUtils::*;
import AXI4Lite_B_Utils::*;
import SpecialRegs::*;
import Cache_Decls::*;
import CacheCorderer::*;
import DReg::*;
import Monitored::*;
import ClientServer::*;
import MemSim::*;
import TieOff::*;
import Fabric_Defs::*;
import StmtFSM::*;
import CPU_IFC::*;
import CHERICap::*;
import CPU_Decode_C::*;
import OneHotArbiter::*;
import CreditCounter::*;
import Bag::*;
import Core_IFC::*;
import AXI4_Common_Types::*;
import GetPut_Aux::*;
import Routable::*;
import SquareRoot::*;
import MemTypesCHERI::*;
import DM_System_Bus::*;
import AXI4_Fake_16550::*;
import TagControllerAXI::*;
import MemBRAM::*;
import Clocks::*;
import SimUtils::*;
import PLIC::*;
import FBox_Core::*;
import MMU_Cache::*;
import CHERICC_Fat::*;
import DM_Common::*;
import SpecialFIFOs::*;
import AXI4_AW_Utils::*;
import MultiLevelTagLookup::*;
import ListExtra::*;
import CPU_Globals::*;
import Debug_Module::*;
import Virtualizable::*;
import FShow::*;
import CSR_MIE::*;
import Assert::*;
import DummyDriver::*;
import Mem::*;
import CPU_Fetch_C::*;
import MasterSlaveCHERI::*;
import Near_Mem_IO_AXI4::*;
import AXI4Lite_W_Utils::*;
import IntMulDiv::*;
import Cur_Cycle::*;
import Semi_FIFOF::*;
import TagTableStructure::*;
import OneWayBus::*;
import TagController::*;
import CSR_RegFile::*;
import FloatingPoint::*;
import MEM::*;
import BRAMCore::*;
import CPU_StageF::*;
import AXI4Lite_Types::*;
import MMU_Cache_Common::*;
import AXI4Lite_Utils::*;
import CSR_RegFile_MSU::*;
import Counter::*;
import AXI4_Types::*;
import AXI4_B_Utils::*;
import ListN::*;
import AXI4Lite_R_Utils::*;
import Cache_Decls_RV64_Sv39_8KB_2way::*;
import FPR_RegFile::*;
import Near_Mem_IFC::*;
import AXI4Stream_Utils::*;
import AXI4Stream::*;

typedef 1 DATASIZE;
typedef 4 ADDRWIDTH;

function Vector #(1, Bool) route_mainBus (r_t x) provisos ( Bits#(r_t,r_l) );
	Bit#(r_l) adress = pack(x);
	Vector#(1, Bool) oneHotAdress = replicate (False);
	// memory -> 0
	if (adress >= 0 && adress < 4096)
		oneHotAdress[0] = True;
	if (adress >= 5096 && adress < 6400)
		oneHotAdress[0] = True;
	return oneHotAdress;
endfunction

module top();
 
	FIFO::FIFO#(Bit#(8)) ff1 <- mkFIFO();
	GetPut::Get#(Bit#(8)) ff1get <- toGet(ff1);
	FIFO::FIFO#(Bit#(8)) ff2 <- mkFIFO();
	GetPut::Put#(Bit#(8)) ff2put <- toPut(ff2);
	Core_IFC::Core_IFC#(SoC_Map::N_External_Interrupt_Sources) core <- mkCore();
	AXI4_Types::AXI4_Slave#(6,64,64,0,0,0,0,0) memory <- mkAXI4SimpleMem(4096, Maybe#("xddd"));

	mkConnection(ff1get,ff2put);
	AXI4_Interconnect::mkAXI4Bus(route_mainBus,mainBus_masters,mainBus_slaves);

endmodule
endpackage
