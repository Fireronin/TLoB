// Example3_tb.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module Example3_tb (
	);

	wire    example3_inst_clk_bfm_clk_clk;       // Example3_inst_clk_bfm:clk -> [Example3_inst:clk_clk, Example3_inst_reset_bfm:clk]
	wire    example3_inst_reset_bfm_reset_reset; // Example3_inst_reset_bfm:reset -> Example3_inst:reset_reset_n

	Example3 example3_inst (
		.clk_clk       (example3_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (example3_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) example3_inst_clk_bfm (
		.clk (example3_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) example3_inst_reset_bfm (
		.reset (example3_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (example3_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
